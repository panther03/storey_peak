// pcie_system.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module pcie_system (
		input  wire        clk_125_clk,                   //          clk_125.clk
		input  wire [31:0] pcie1_hip_ctrl_test_in,        //   pcie1_hip_ctrl.test_in
		input  wire        pcie1_hip_ctrl_simu_mode_pipe, //                 .simu_mode_pipe
		input  wire        pcie1_hip_serial_rx_in0,       // pcie1_hip_serial.rx_in0
		input  wire        pcie1_hip_serial_rx_in1,       //                 .rx_in1
		input  wire        pcie1_hip_serial_rx_in2,       //                 .rx_in2
		input  wire        pcie1_hip_serial_rx_in3,       //                 .rx_in3
		input  wire        pcie1_hip_serial_rx_in4,       //                 .rx_in4
		input  wire        pcie1_hip_serial_rx_in5,       //                 .rx_in5
		input  wire        pcie1_hip_serial_rx_in6,       //                 .rx_in6
		input  wire        pcie1_hip_serial_rx_in7,       //                 .rx_in7
		output wire        pcie1_hip_serial_tx_out0,      //                 .tx_out0
		output wire        pcie1_hip_serial_tx_out1,      //                 .tx_out1
		output wire        pcie1_hip_serial_tx_out2,      //                 .tx_out2
		output wire        pcie1_hip_serial_tx_out3,      //                 .tx_out3
		output wire        pcie1_hip_serial_tx_out4,      //                 .tx_out4
		output wire        pcie1_hip_serial_tx_out5,      //                 .tx_out5
		output wire        pcie1_hip_serial_tx_out6,      //                 .tx_out6
		output wire        pcie1_hip_serial_tx_out7,      //                 .tx_out7
		input  wire        pcie1_npor_npor,               //       pcie1_npor.npor
		input  wire        pcie1_npor_pin_perst,          //                 .pin_perst
		input  wire        pcie1_refclk_clk,              //     pcie1_refclk.clk
		input  wire [31:0] pcie2_hip_ctrl_test_in,        //   pcie2_hip_ctrl.test_in
		input  wire        pcie2_hip_ctrl_simu_mode_pipe, //                 .simu_mode_pipe
		input  wire        pcie2_hip_serial_rx_in0,       // pcie2_hip_serial.rx_in0
		input  wire        pcie2_hip_serial_rx_in1,       //                 .rx_in1
		input  wire        pcie2_hip_serial_rx_in2,       //                 .rx_in2
		input  wire        pcie2_hip_serial_rx_in3,       //                 .rx_in3
		input  wire        pcie2_hip_serial_rx_in4,       //                 .rx_in4
		input  wire        pcie2_hip_serial_rx_in5,       //                 .rx_in5
		input  wire        pcie2_hip_serial_rx_in6,       //                 .rx_in6
		input  wire        pcie2_hip_serial_rx_in7,       //                 .rx_in7
		output wire        pcie2_hip_serial_tx_out0,      //                 .tx_out0
		output wire        pcie2_hip_serial_tx_out1,      //                 .tx_out1
		output wire        pcie2_hip_serial_tx_out2,      //                 .tx_out2
		output wire        pcie2_hip_serial_tx_out3,      //                 .tx_out3
		output wire        pcie2_hip_serial_tx_out4,      //                 .tx_out4
		output wire        pcie2_hip_serial_tx_out5,      //                 .tx_out5
		output wire        pcie2_hip_serial_tx_out6,      //                 .tx_out6
		output wire        pcie2_hip_serial_tx_out7,      //                 .tx_out7
		input  wire        pcie2_npor_npor,               //       pcie2_npor.npor
		input  wire        pcie2_npor_pin_perst,          //                 .pin_perst
		input  wire        pcie2_refclk_clk,              //     pcie2_refclk.clk
		input  wire        rst_125_reset_n,               //          rst_125.reset_n
		input  wire        uart_conduit_rxd,              //     uart_conduit.rxd
		output wire        uart_conduit_txd               //                 .txd
	);

	wire          pcie1_coreclkout_clk;                                  // pcie1:coreclkout -> [intel_lw_uart_0:clk, mm_interconnect_0:pcie1_coreclkout_clk, rst_controller_001:clk, rst_controller_002:clk, sysid_qsys_0:clock]
	wire  [459:0] pcie2_reconfig_from_xcvr_reconfig_from_xcvr;           // pcie2:reconfig_from_xcvr -> alt_xcvr_reconfig_1:reconfig_from_xcvr
	wire  [459:0] pcie1_reconfig_from_xcvr_reconfig_from_xcvr;           // pcie1:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [699:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr; // alt_xcvr_reconfig_0:reconfig_to_xcvr -> pcie1:reconfig_to_xcvr
	wire  [699:0] alt_xcvr_reconfig_1_reconfig_to_xcvr_reconfig_to_xcvr; // alt_xcvr_reconfig_1:reconfig_to_xcvr -> pcie2:reconfig_to_xcvr
	wire          pcie1_rxm_bar0_waitrequest;                            // mm_interconnect_0:pcie1_Rxm_BAR0_waitrequest -> pcie1:RxmWaitRequest_0_i
	wire  [127:0] pcie1_rxm_bar0_readdata;                               // mm_interconnect_0:pcie1_Rxm_BAR0_readdata -> pcie1:RxmReadData_0_i
	wire   [31:0] pcie1_rxm_bar0_address;                                // pcie1:RxmAddress_0_o -> mm_interconnect_0:pcie1_Rxm_BAR0_address
	wire          pcie1_rxm_bar0_read;                                   // pcie1:RxmRead_0_o -> mm_interconnect_0:pcie1_Rxm_BAR0_read
	wire   [15:0] pcie1_rxm_bar0_byteenable;                             // pcie1:RxmByteEnable_0_o -> mm_interconnect_0:pcie1_Rxm_BAR0_byteenable
	wire          pcie1_rxm_bar0_readdatavalid;                          // mm_interconnect_0:pcie1_Rxm_BAR0_readdatavalid -> pcie1:RxmReadDataValid_0_i
	wire          pcie1_rxm_bar0_write;                                  // pcie1:RxmWrite_0_o -> mm_interconnect_0:pcie1_Rxm_BAR0_write
	wire  [127:0] pcie1_rxm_bar0_writedata;                              // pcie1:RxmWriteData_0_o -> mm_interconnect_0:pcie1_Rxm_BAR0_writedata
	wire    [5:0] pcie1_rxm_bar0_burstcount;                             // pcie1:RxmBurstCount_0_o -> mm_interconnect_0:pcie1_Rxm_BAR0_burstcount
	wire   [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [15:0] mm_interconnect_0_intel_lw_uart_0_s1_readdata;         // intel_lw_uart_0:readdata -> mm_interconnect_0:intel_lw_uart_0_s1_readdata
	wire    [2:0] mm_interconnect_0_intel_lw_uart_0_s1_address;          // mm_interconnect_0:intel_lw_uart_0_s1_address -> intel_lw_uart_0:address
	wire          mm_interconnect_0_intel_lw_uart_0_s1_read;             // mm_interconnect_0:intel_lw_uart_0_s1_read -> intel_lw_uart_0:read
	wire          mm_interconnect_0_intel_lw_uart_0_s1_write;            // mm_interconnect_0:intel_lw_uart_0_s1_write -> intel_lw_uart_0:write
	wire   [15:0] mm_interconnect_0_intel_lw_uart_0_s1_writedata;        // mm_interconnect_0:intel_lw_uart_0_s1_writedata -> intel_lw_uart_0:writedata
	wire          rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, alt_xcvr_reconfig_1:mgmt_rst_reset]
	wire          rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> [intel_lw_uart_0:reset_n, mm_interconnect_0:intel_lw_uart_0_reset_reset_bridge_in_reset_reset]
	wire          pcie1_nreset_status_reset;                             // pcie1:reset_status -> [rst_controller_001:reset_in0, rst_controller_002:reset_in1]
	wire          rst_controller_002_reset_out_reset;                    // rst_controller_002:reset_out -> [mm_interconnect_0:sysid_qsys_0_reset_reset_bridge_in_reset_reset, sysid_qsys_0:reset_n]

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (10),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (),                                                      //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_125_clk),                                           //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                        //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (),                                                      //      reconfig_mgmt.address
		.reconfig_mgmt_read        (),                                                      //                   .read
		.reconfig_mgmt_readdata    (),                                                      //                   .readdata
		.reconfig_mgmt_waitrequest (),                                                      //                   .waitrequest
		.reconfig_mgmt_write       (),                                                      //                   .write
		.reconfig_mgmt_writedata   (),                                                      //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie1_reconfig_from_xcvr_reconfig_from_xcvr),           // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                      //        (terminated)
		.rx_cal_busy               (),                                                      //        (terminated)
		.cal_busy_in               (1'b0),                                                  //        (terminated)
		.reconfig_mif_address      (),                                                      //        (terminated)
		.reconfig_mif_read         (),                                                      //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                  //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                   //        (terminated)
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (10),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_1 (
		.reconfig_busy             (),                                                      //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_125_clk),                                           //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                        //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (),                                                      //      reconfig_mgmt.address
		.reconfig_mgmt_read        (),                                                      //                   .read
		.reconfig_mgmt_readdata    (),                                                      //                   .readdata
		.reconfig_mgmt_waitrequest (),                                                      //                   .waitrequest
		.reconfig_mgmt_write       (),                                                      //                   .write
		.reconfig_mgmt_writedata   (),                                                      //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_1_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie2_reconfig_from_xcvr_reconfig_from_xcvr),           // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                      //        (terminated)
		.rx_cal_busy               (),                                                      //        (terminated)
		.cal_busy_in               (1'b0),                                                  //        (terminated)
		.reconfig_mif_address      (),                                                      //        (terminated)
		.reconfig_mif_read         (),                                                      //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                  //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                   //        (terminated)
	);

	intel_lw_uart #(
		.dataBits                     (8),
		.fixedBaud                    (1),
		.parity                       ("NONE"),
		.stopBits                     (1),
		.syncRegDepth                 (2),
		.useCtsRts                    (0),
		.useEopRegister               (0),
		.useRegTXFIFO                 (0),
		.useRegRXFIFO                 (0),
		.simTrueBaud                  (0),
		.divisorConstant              (2169),
		.divisorConstantWidth         (12),
		.derivedTxfifoDepth           (2048),
		.derivedRxfifoDepth           (2048),
		.derivedRxfifoAlmostFullValue (2047),
		.txfifoWidthu                 (11),
		.rxfifoWidthu                 (11)
	) intel_lw_uart_0 (
		.clk       (pcie1_coreclkout_clk),                           //                 clk.clk
		.reset_n   (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address   (mm_interconnect_0_intel_lw_uart_0_s1_address),   //                  s1.address
		.read      (mm_interconnect_0_intel_lw_uart_0_s1_read),      //                    .read
		.write     (mm_interconnect_0_intel_lw_uart_0_s1_write),     //                    .write
		.writedata (mm_interconnect_0_intel_lw_uart_0_s1_writedata), //                    .writedata
		.readdata  (mm_interconnect_0_intel_lw_uart_0_s1_readdata),  //                    .readdata
		.rxd       (uart_conduit_rxd),                               // external_connection.rxd
		.txd       (uart_conduit_txd),                               //                    .txd
		.irq       (),                                               //                 irq.irq
		.cts_n     (1'b1),                                           //         (terminated)
		.rts_n     ()                                                //         (terminated)
	);

	altpcie_sv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen2 (5.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.enable_power_on_rst_pulse_hwtcl          (0),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (6),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (0),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (167),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (418),
		.subsystem_device_id_hwtcl                (1),
		.max_payload_size_hwtcl                   (128),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (4466),
		.vsec_rev_hwtcl                           (0),
		.user_id_hwtcl                            (0),
		.avmm_width_hwtcl                         (128),
		.AVALON_ADDR_WIDTH                        (32),
		.avmm_burst_width_hwtcl                   (6),
		.CB_PCIE_MODE                             (1),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (128),
		.CG_AVALON_S_ADDR_WIDTH                   (21),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (0),
		.CG_ENABLE_ADVANCED_INTERRUPT             (0),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (2),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (20),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (248500),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.hip_reconfig_hwtcl                       (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (700),
		.reconfig_from_xcvr_width                 (460),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (0),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15)
	) pcie1 (
		.coreclkout           (pcie1_coreclkout_clk),                                  //          coreclkout.clk
		.refclk               (pcie1_refclk_clk),                                      //              refclk.clk
		.npor                 (pcie1_npor_npor),                                       //                npor.npor
		.pin_perst            (pcie1_npor_pin_perst),                                  //                    .pin_perst
		.reset_status         (pcie1_nreset_status_reset),                             //       nreset_status.reset_n
		.RxmAddress_0_o       (pcie1_rxm_bar0_address),                                //            Rxm_BAR0.address
		.RxmRead_0_o          (pcie1_rxm_bar0_read),                                   //                    .read
		.RxmWaitRequest_0_i   (pcie1_rxm_bar0_waitrequest),                            //                    .waitrequest
		.RxmWrite_0_o         (pcie1_rxm_bar0_write),                                  //                    .write
		.RxmReadDataValid_0_i (pcie1_rxm_bar0_readdatavalid),                          //                    .readdatavalid
		.RxmReadData_0_i      (pcie1_rxm_bar0_readdata),                               //                    .readdata
		.RxmWriteData_0_o     (pcie1_rxm_bar0_writedata),                              //                    .writedata
		.RxmBurstCount_0_o    (pcie1_rxm_bar0_burstcount),                             //                    .burstcount
		.RxmByteEnable_0_o    (pcie1_rxm_bar0_byteenable),                             //                    .byteenable
		.derr_cor_ext_rcv     (),                                                      //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (),                                                      //                    .derr_cor_ext_rpl
		.derr_rpl             (),                                                      //                    .derr_rpl
		.dlup                 (),                                                      //                    .dlup
		.dlup_exit            (),                                                      //                    .dlup_exit
		.ev128ns              (),                                                      //                    .ev128ns
		.ev1us                (),                                                      //                    .ev1us
		.hotrst_exit          (),                                                      //                    .hotrst_exit
		.int_status           (),                                                      //                    .int_status
		.l2_exit              (),                                                      //                    .l2_exit
		.lane_act             (),                                                      //                    .lane_act
		.ltssmstate           (),                                                      //                    .ltssmstate
		.rx_par_err           (),                                                      //                    .rx_par_err
		.tx_par_err           (),                                                      //                    .tx_par_err
		.cfg_par_err          (),                                                      //                    .cfg_par_err
		.ko_cpl_spc_header    (),                                                      //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (),                                                      //                    .ko_cpl_spc_data
		.currentspeed         (),                                                      //    hip_currentspeed.currentspeed
		.reconfig_to_xcvr     (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (pcie1_reconfig_from_xcvr_reconfig_from_xcvr),           //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (),                                                      // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (pcie1_hip_serial_rx_in0),                               //          hip_serial.rx_in0
		.rx_in1               (pcie1_hip_serial_rx_in1),                               //                    .rx_in1
		.rx_in2               (pcie1_hip_serial_rx_in2),                               //                    .rx_in2
		.rx_in3               (pcie1_hip_serial_rx_in3),                               //                    .rx_in3
		.rx_in4               (pcie1_hip_serial_rx_in4),                               //                    .rx_in4
		.rx_in5               (pcie1_hip_serial_rx_in5),                               //                    .rx_in5
		.rx_in6               (pcie1_hip_serial_rx_in6),                               //                    .rx_in6
		.rx_in7               (pcie1_hip_serial_rx_in7),                               //                    .rx_in7
		.tx_out0              (pcie1_hip_serial_tx_out0),                              //                    .tx_out0
		.tx_out1              (pcie1_hip_serial_tx_out1),                              //                    .tx_out1
		.tx_out2              (pcie1_hip_serial_tx_out2),                              //                    .tx_out2
		.tx_out3              (pcie1_hip_serial_tx_out3),                              //                    .tx_out3
		.tx_out4              (pcie1_hip_serial_tx_out4),                              //                    .tx_out4
		.tx_out5              (pcie1_hip_serial_tx_out5),                              //                    .tx_out5
		.tx_out6              (pcie1_hip_serial_tx_out6),                              //                    .tx_out6
		.tx_out7              (pcie1_hip_serial_tx_out7),                              //                    .tx_out7
		.sim_pipe_pclk_in     (),                                                      //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                                      //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                                      //                    .sim_ltssmstate
		.eidleinfersel0       (),                                                      //                    .eidleinfersel0
		.eidleinfersel1       (),                                                      //                    .eidleinfersel1
		.eidleinfersel2       (),                                                      //                    .eidleinfersel2
		.eidleinfersel3       (),                                                      //                    .eidleinfersel3
		.eidleinfersel4       (),                                                      //                    .eidleinfersel4
		.eidleinfersel5       (),                                                      //                    .eidleinfersel5
		.eidleinfersel6       (),                                                      //                    .eidleinfersel6
		.eidleinfersel7       (),                                                      //                    .eidleinfersel7
		.powerdown0           (),                                                      //                    .powerdown0
		.powerdown1           (),                                                      //                    .powerdown1
		.powerdown2           (),                                                      //                    .powerdown2
		.powerdown3           (),                                                      //                    .powerdown3
		.powerdown4           (),                                                      //                    .powerdown4
		.powerdown5           (),                                                      //                    .powerdown5
		.powerdown6           (),                                                      //                    .powerdown6
		.powerdown7           (),                                                      //                    .powerdown7
		.rxpolarity0          (),                                                      //                    .rxpolarity0
		.rxpolarity1          (),                                                      //                    .rxpolarity1
		.rxpolarity2          (),                                                      //                    .rxpolarity2
		.rxpolarity3          (),                                                      //                    .rxpolarity3
		.rxpolarity4          (),                                                      //                    .rxpolarity4
		.rxpolarity5          (),                                                      //                    .rxpolarity5
		.rxpolarity6          (),                                                      //                    .rxpolarity6
		.rxpolarity7          (),                                                      //                    .rxpolarity7
		.txcompl0             (),                                                      //                    .txcompl0
		.txcompl1             (),                                                      //                    .txcompl1
		.txcompl2             (),                                                      //                    .txcompl2
		.txcompl3             (),                                                      //                    .txcompl3
		.txcompl4             (),                                                      //                    .txcompl4
		.txcompl5             (),                                                      //                    .txcompl5
		.txcompl6             (),                                                      //                    .txcompl6
		.txcompl7             (),                                                      //                    .txcompl7
		.txdata0              (),                                                      //                    .txdata0
		.txdata1              (),                                                      //                    .txdata1
		.txdata2              (),                                                      //                    .txdata2
		.txdata3              (),                                                      //                    .txdata3
		.txdata4              (),                                                      //                    .txdata4
		.txdata5              (),                                                      //                    .txdata5
		.txdata6              (),                                                      //                    .txdata6
		.txdata7              (),                                                      //                    .txdata7
		.txdatak0             (),                                                      //                    .txdatak0
		.txdatak1             (),                                                      //                    .txdatak1
		.txdatak2             (),                                                      //                    .txdatak2
		.txdatak3             (),                                                      //                    .txdatak3
		.txdatak4             (),                                                      //                    .txdatak4
		.txdatak5             (),                                                      //                    .txdatak5
		.txdatak6             (),                                                      //                    .txdatak6
		.txdatak7             (),                                                      //                    .txdatak7
		.txdetectrx0          (),                                                      //                    .txdetectrx0
		.txdetectrx1          (),                                                      //                    .txdetectrx1
		.txdetectrx2          (),                                                      //                    .txdetectrx2
		.txdetectrx3          (),                                                      //                    .txdetectrx3
		.txdetectrx4          (),                                                      //                    .txdetectrx4
		.txdetectrx5          (),                                                      //                    .txdetectrx5
		.txdetectrx6          (),                                                      //                    .txdetectrx6
		.txdetectrx7          (),                                                      //                    .txdetectrx7
		.txelecidle0          (),                                                      //                    .txelecidle0
		.txelecidle1          (),                                                      //                    .txelecidle1
		.txelecidle2          (),                                                      //                    .txelecidle2
		.txelecidle3          (),                                                      //                    .txelecidle3
		.txelecidle4          (),                                                      //                    .txelecidle4
		.txelecidle5          (),                                                      //                    .txelecidle5
		.txelecidle6          (),                                                      //                    .txelecidle6
		.txelecidle7          (),                                                      //                    .txelecidle7
		.txdeemph0            (),                                                      //                    .txdeemph0
		.txdeemph1            (),                                                      //                    .txdeemph1
		.txdeemph2            (),                                                      //                    .txdeemph2
		.txdeemph3            (),                                                      //                    .txdeemph3
		.txdeemph4            (),                                                      //                    .txdeemph4
		.txdeemph5            (),                                                      //                    .txdeemph5
		.txdeemph6            (),                                                      //                    .txdeemph6
		.txdeemph7            (),                                                      //                    .txdeemph7
		.txmargin0            (),                                                      //                    .txmargin0
		.txmargin1            (),                                                      //                    .txmargin1
		.txmargin2            (),                                                      //                    .txmargin2
		.txmargin3            (),                                                      //                    .txmargin3
		.txmargin4            (),                                                      //                    .txmargin4
		.txmargin5            (),                                                      //                    .txmargin5
		.txmargin6            (),                                                      //                    .txmargin6
		.txmargin7            (),                                                      //                    .txmargin7
		.txswing0             (),                                                      //                    .txswing0
		.txswing1             (),                                                      //                    .txswing1
		.txswing2             (),                                                      //                    .txswing2
		.txswing3             (),                                                      //                    .txswing3
		.txswing4             (),                                                      //                    .txswing4
		.txswing5             (),                                                      //                    .txswing5
		.txswing6             (),                                                      //                    .txswing6
		.txswing7             (),                                                      //                    .txswing7
		.phystatus0           (),                                                      //                    .phystatus0
		.phystatus1           (),                                                      //                    .phystatus1
		.phystatus2           (),                                                      //                    .phystatus2
		.phystatus3           (),                                                      //                    .phystatus3
		.phystatus4           (),                                                      //                    .phystatus4
		.phystatus5           (),                                                      //                    .phystatus5
		.phystatus6           (),                                                      //                    .phystatus6
		.phystatus7           (),                                                      //                    .phystatus7
		.rxdata0              (),                                                      //                    .rxdata0
		.rxdata1              (),                                                      //                    .rxdata1
		.rxdata2              (),                                                      //                    .rxdata2
		.rxdata3              (),                                                      //                    .rxdata3
		.rxdata4              (),                                                      //                    .rxdata4
		.rxdata5              (),                                                      //                    .rxdata5
		.rxdata6              (),                                                      //                    .rxdata6
		.rxdata7              (),                                                      //                    .rxdata7
		.rxdatak0             (),                                                      //                    .rxdatak0
		.rxdatak1             (),                                                      //                    .rxdatak1
		.rxdatak2             (),                                                      //                    .rxdatak2
		.rxdatak3             (),                                                      //                    .rxdatak3
		.rxdatak4             (),                                                      //                    .rxdatak4
		.rxdatak5             (),                                                      //                    .rxdatak5
		.rxdatak6             (),                                                      //                    .rxdatak6
		.rxdatak7             (),                                                      //                    .rxdatak7
		.rxelecidle0          (),                                                      //                    .rxelecidle0
		.rxelecidle1          (),                                                      //                    .rxelecidle1
		.rxelecidle2          (),                                                      //                    .rxelecidle2
		.rxelecidle3          (),                                                      //                    .rxelecidle3
		.rxelecidle4          (),                                                      //                    .rxelecidle4
		.rxelecidle5          (),                                                      //                    .rxelecidle5
		.rxelecidle6          (),                                                      //                    .rxelecidle6
		.rxelecidle7          (),                                                      //                    .rxelecidle7
		.rxstatus0            (),                                                      //                    .rxstatus0
		.rxstatus1            (),                                                      //                    .rxstatus1
		.rxstatus2            (),                                                      //                    .rxstatus2
		.rxstatus3            (),                                                      //                    .rxstatus3
		.rxstatus4            (),                                                      //                    .rxstatus4
		.rxstatus5            (),                                                      //                    .rxstatus5
		.rxstatus6            (),                                                      //                    .rxstatus6
		.rxstatus7            (),                                                      //                    .rxstatus7
		.rxvalid0             (),                                                      //                    .rxvalid0
		.rxvalid1             (),                                                      //                    .rxvalid1
		.rxvalid2             (),                                                      //                    .rxvalid2
		.rxvalid3             (),                                                      //                    .rxvalid3
		.rxvalid4             (),                                                      //                    .rxvalid4
		.rxvalid5             (),                                                      //                    .rxvalid5
		.rxvalid6             (),                                                      //                    .rxvalid6
		.rxvalid7             (),                                                      //                    .rxvalid7
		.test_in              (pcie1_hip_ctrl_test_in),                                //            hip_ctrl.test_in
		.simu_mode_pipe       (pcie1_hip_ctrl_simu_mode_pipe),                         //                    .simu_mode_pipe
		.rxdataskip0          (1'b0),                                                  //         (terminated)
		.rxdataskip1          (1'b0),                                                  //         (terminated)
		.rxdataskip2          (1'b0),                                                  //         (terminated)
		.rxdataskip3          (1'b0),                                                  //         (terminated)
		.rxdataskip4          (1'b0),                                                  //         (terminated)
		.rxdataskip5          (1'b0),                                                  //         (terminated)
		.rxdataskip6          (1'b0),                                                  //         (terminated)
		.rxdataskip7          (1'b0),                                                  //         (terminated)
		.rxblkst0             (1'b0),                                                  //         (terminated)
		.rxblkst1             (1'b0),                                                  //         (terminated)
		.rxblkst2             (1'b0),                                                  //         (terminated)
		.rxblkst3             (1'b0),                                                  //         (terminated)
		.rxblkst4             (1'b0),                                                  //         (terminated)
		.rxblkst5             (1'b0),                                                  //         (terminated)
		.rxblkst6             (1'b0),                                                  //         (terminated)
		.rxblkst7             (1'b0),                                                  //         (terminated)
		.rxsynchd0            (2'b00),                                                 //         (terminated)
		.rxsynchd1            (2'b00),                                                 //         (terminated)
		.rxsynchd2            (2'b00),                                                 //         (terminated)
		.rxsynchd3            (2'b00),                                                 //         (terminated)
		.rxsynchd4            (2'b00),                                                 //         (terminated)
		.rxsynchd5            (2'b00),                                                 //         (terminated)
		.rxsynchd6            (2'b00),                                                 //         (terminated)
		.rxsynchd7            (2'b00),                                                 //         (terminated)
		.rxfreqlocked0        (1'b0),                                                  //         (terminated)
		.rxfreqlocked1        (1'b0),                                                  //         (terminated)
		.rxfreqlocked2        (1'b0),                                                  //         (terminated)
		.rxfreqlocked3        (1'b0),                                                  //         (terminated)
		.rxfreqlocked4        (1'b0),                                                  //         (terminated)
		.rxfreqlocked5        (1'b0),                                                  //         (terminated)
		.rxfreqlocked6        (1'b0),                                                  //         (terminated)
		.rxfreqlocked7        (1'b0),                                                  //         (terminated)
		.currentcoeff0        (),                                                      //         (terminated)
		.currentcoeff1        (),                                                      //         (terminated)
		.currentcoeff2        (),                                                      //         (terminated)
		.currentcoeff3        (),                                                      //         (terminated)
		.currentcoeff4        (),                                                      //         (terminated)
		.currentcoeff5        (),                                                      //         (terminated)
		.currentcoeff6        (),                                                      //         (terminated)
		.currentcoeff7        (),                                                      //         (terminated)
		.currentrxpreset0     (),                                                      //         (terminated)
		.currentrxpreset1     (),                                                      //         (terminated)
		.currentrxpreset2     (),                                                      //         (terminated)
		.currentrxpreset3     (),                                                      //         (terminated)
		.currentrxpreset4     (),                                                      //         (terminated)
		.currentrxpreset5     (),                                                      //         (terminated)
		.currentrxpreset6     (),                                                      //         (terminated)
		.currentrxpreset7     (),                                                      //         (terminated)
		.txsynchd0            (),                                                      //         (terminated)
		.txsynchd1            (),                                                      //         (terminated)
		.txsynchd2            (),                                                      //         (terminated)
		.txsynchd3            (),                                                      //         (terminated)
		.txsynchd4            (),                                                      //         (terminated)
		.txsynchd5            (),                                                      //         (terminated)
		.txsynchd6            (),                                                      //         (terminated)
		.txsynchd7            (),                                                      //         (terminated)
		.txblkst0             (),                                                      //         (terminated)
		.txblkst1             (),                                                      //         (terminated)
		.txblkst2             (),                                                      //         (terminated)
		.txblkst3             (),                                                      //         (terminated)
		.txblkst4             (),                                                      //         (terminated)
		.txblkst5             (),                                                      //         (terminated)
		.txblkst6             (),                                                      //         (terminated)
		.txblkst7             ()                                                       //         (terminated)
	);

	altpcie_sv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen2 (5.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.enable_power_on_rst_pulse_hwtcl          (0),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (0),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (0),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (167),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (418),
		.subsystem_device_id_hwtcl                (0),
		.max_payload_size_hwtcl                   (128),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (4466),
		.vsec_rev_hwtcl                           (0),
		.user_id_hwtcl                            (0),
		.avmm_width_hwtcl                         (128),
		.AVALON_ADDR_WIDTH                        (32),
		.avmm_burst_width_hwtcl                   (6),
		.CB_PCIE_MODE                             (1),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (128),
		.CG_AVALON_S_ADDR_WIDTH                   (21),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (0),
		.CG_ENABLE_ADVANCED_INTERRUPT             (0),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (2),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (20),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (248500),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.hip_reconfig_hwtcl                       (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (700),
		.reconfig_from_xcvr_width                 (460),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (0),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15)
	) pcie2 (
		.coreclkout           (),                                                      //          coreclkout.clk
		.refclk               (pcie2_refclk_clk),                                      //              refclk.clk
		.npor                 (pcie2_npor_npor),                                       //                npor.npor
		.pin_perst            (pcie2_npor_pin_perst),                                  //                    .pin_perst
		.reset_status         (),                                                      //       nreset_status.reset_n
		.RxmAddress_0_o       (),                                                      //            Rxm_BAR0.address
		.RxmRead_0_o          (),                                                      //                    .read
		.RxmWaitRequest_0_i   (),                                                      //                    .waitrequest
		.RxmWrite_0_o         (),                                                      //                    .write
		.RxmReadDataValid_0_i (),                                                      //                    .readdatavalid
		.RxmReadData_0_i      (),                                                      //                    .readdata
		.RxmWriteData_0_o     (),                                                      //                    .writedata
		.RxmBurstCount_0_o    (),                                                      //                    .burstcount
		.RxmByteEnable_0_o    (),                                                      //                    .byteenable
		.derr_cor_ext_rcv     (),                                                      //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (),                                                      //                    .derr_cor_ext_rpl
		.derr_rpl             (),                                                      //                    .derr_rpl
		.dlup                 (),                                                      //                    .dlup
		.dlup_exit            (),                                                      //                    .dlup_exit
		.ev128ns              (),                                                      //                    .ev128ns
		.ev1us                (),                                                      //                    .ev1us
		.hotrst_exit          (),                                                      //                    .hotrst_exit
		.int_status           (),                                                      //                    .int_status
		.l2_exit              (),                                                      //                    .l2_exit
		.lane_act             (),                                                      //                    .lane_act
		.ltssmstate           (),                                                      //                    .ltssmstate
		.rx_par_err           (),                                                      //                    .rx_par_err
		.tx_par_err           (),                                                      //                    .tx_par_err
		.cfg_par_err          (),                                                      //                    .cfg_par_err
		.ko_cpl_spc_header    (),                                                      //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (),                                                      //                    .ko_cpl_spc_data
		.currentspeed         (),                                                      //    hip_currentspeed.currentspeed
		.reconfig_to_xcvr     (alt_xcvr_reconfig_1_reconfig_to_xcvr_reconfig_to_xcvr), //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (pcie2_reconfig_from_xcvr_reconfig_from_xcvr),           //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (),                                                      // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (pcie2_hip_serial_rx_in0),                               //          hip_serial.rx_in0
		.rx_in1               (pcie2_hip_serial_rx_in1),                               //                    .rx_in1
		.rx_in2               (pcie2_hip_serial_rx_in2),                               //                    .rx_in2
		.rx_in3               (pcie2_hip_serial_rx_in3),                               //                    .rx_in3
		.rx_in4               (pcie2_hip_serial_rx_in4),                               //                    .rx_in4
		.rx_in5               (pcie2_hip_serial_rx_in5),                               //                    .rx_in5
		.rx_in6               (pcie2_hip_serial_rx_in6),                               //                    .rx_in6
		.rx_in7               (pcie2_hip_serial_rx_in7),                               //                    .rx_in7
		.tx_out0              (pcie2_hip_serial_tx_out0),                              //                    .tx_out0
		.tx_out1              (pcie2_hip_serial_tx_out1),                              //                    .tx_out1
		.tx_out2              (pcie2_hip_serial_tx_out2),                              //                    .tx_out2
		.tx_out3              (pcie2_hip_serial_tx_out3),                              //                    .tx_out3
		.tx_out4              (pcie2_hip_serial_tx_out4),                              //                    .tx_out4
		.tx_out5              (pcie2_hip_serial_tx_out5),                              //                    .tx_out5
		.tx_out6              (pcie2_hip_serial_tx_out6),                              //                    .tx_out6
		.tx_out7              (pcie2_hip_serial_tx_out7),                              //                    .tx_out7
		.sim_pipe_pclk_in     (),                                                      //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                                      //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                                      //                    .sim_ltssmstate
		.eidleinfersel0       (),                                                      //                    .eidleinfersel0
		.eidleinfersel1       (),                                                      //                    .eidleinfersel1
		.eidleinfersel2       (),                                                      //                    .eidleinfersel2
		.eidleinfersel3       (),                                                      //                    .eidleinfersel3
		.eidleinfersel4       (),                                                      //                    .eidleinfersel4
		.eidleinfersel5       (),                                                      //                    .eidleinfersel5
		.eidleinfersel6       (),                                                      //                    .eidleinfersel6
		.eidleinfersel7       (),                                                      //                    .eidleinfersel7
		.powerdown0           (),                                                      //                    .powerdown0
		.powerdown1           (),                                                      //                    .powerdown1
		.powerdown2           (),                                                      //                    .powerdown2
		.powerdown3           (),                                                      //                    .powerdown3
		.powerdown4           (),                                                      //                    .powerdown4
		.powerdown5           (),                                                      //                    .powerdown5
		.powerdown6           (),                                                      //                    .powerdown6
		.powerdown7           (),                                                      //                    .powerdown7
		.rxpolarity0          (),                                                      //                    .rxpolarity0
		.rxpolarity1          (),                                                      //                    .rxpolarity1
		.rxpolarity2          (),                                                      //                    .rxpolarity2
		.rxpolarity3          (),                                                      //                    .rxpolarity3
		.rxpolarity4          (),                                                      //                    .rxpolarity4
		.rxpolarity5          (),                                                      //                    .rxpolarity5
		.rxpolarity6          (),                                                      //                    .rxpolarity6
		.rxpolarity7          (),                                                      //                    .rxpolarity7
		.txcompl0             (),                                                      //                    .txcompl0
		.txcompl1             (),                                                      //                    .txcompl1
		.txcompl2             (),                                                      //                    .txcompl2
		.txcompl3             (),                                                      //                    .txcompl3
		.txcompl4             (),                                                      //                    .txcompl4
		.txcompl5             (),                                                      //                    .txcompl5
		.txcompl6             (),                                                      //                    .txcompl6
		.txcompl7             (),                                                      //                    .txcompl7
		.txdata0              (),                                                      //                    .txdata0
		.txdata1              (),                                                      //                    .txdata1
		.txdata2              (),                                                      //                    .txdata2
		.txdata3              (),                                                      //                    .txdata3
		.txdata4              (),                                                      //                    .txdata4
		.txdata5              (),                                                      //                    .txdata5
		.txdata6              (),                                                      //                    .txdata6
		.txdata7              (),                                                      //                    .txdata7
		.txdatak0             (),                                                      //                    .txdatak0
		.txdatak1             (),                                                      //                    .txdatak1
		.txdatak2             (),                                                      //                    .txdatak2
		.txdatak3             (),                                                      //                    .txdatak3
		.txdatak4             (),                                                      //                    .txdatak4
		.txdatak5             (),                                                      //                    .txdatak5
		.txdatak6             (),                                                      //                    .txdatak6
		.txdatak7             (),                                                      //                    .txdatak7
		.txdetectrx0          (),                                                      //                    .txdetectrx0
		.txdetectrx1          (),                                                      //                    .txdetectrx1
		.txdetectrx2          (),                                                      //                    .txdetectrx2
		.txdetectrx3          (),                                                      //                    .txdetectrx3
		.txdetectrx4          (),                                                      //                    .txdetectrx4
		.txdetectrx5          (),                                                      //                    .txdetectrx5
		.txdetectrx6          (),                                                      //                    .txdetectrx6
		.txdetectrx7          (),                                                      //                    .txdetectrx7
		.txelecidle0          (),                                                      //                    .txelecidle0
		.txelecidle1          (),                                                      //                    .txelecidle1
		.txelecidle2          (),                                                      //                    .txelecidle2
		.txelecidle3          (),                                                      //                    .txelecidle3
		.txelecidle4          (),                                                      //                    .txelecidle4
		.txelecidle5          (),                                                      //                    .txelecidle5
		.txelecidle6          (),                                                      //                    .txelecidle6
		.txelecidle7          (),                                                      //                    .txelecidle7
		.txdeemph0            (),                                                      //                    .txdeemph0
		.txdeemph1            (),                                                      //                    .txdeemph1
		.txdeemph2            (),                                                      //                    .txdeemph2
		.txdeemph3            (),                                                      //                    .txdeemph3
		.txdeemph4            (),                                                      //                    .txdeemph4
		.txdeemph5            (),                                                      //                    .txdeemph5
		.txdeemph6            (),                                                      //                    .txdeemph6
		.txdeemph7            (),                                                      //                    .txdeemph7
		.txmargin0            (),                                                      //                    .txmargin0
		.txmargin1            (),                                                      //                    .txmargin1
		.txmargin2            (),                                                      //                    .txmargin2
		.txmargin3            (),                                                      //                    .txmargin3
		.txmargin4            (),                                                      //                    .txmargin4
		.txmargin5            (),                                                      //                    .txmargin5
		.txmargin6            (),                                                      //                    .txmargin6
		.txmargin7            (),                                                      //                    .txmargin7
		.txswing0             (),                                                      //                    .txswing0
		.txswing1             (),                                                      //                    .txswing1
		.txswing2             (),                                                      //                    .txswing2
		.txswing3             (),                                                      //                    .txswing3
		.txswing4             (),                                                      //                    .txswing4
		.txswing5             (),                                                      //                    .txswing5
		.txswing6             (),                                                      //                    .txswing6
		.txswing7             (),                                                      //                    .txswing7
		.phystatus0           (),                                                      //                    .phystatus0
		.phystatus1           (),                                                      //                    .phystatus1
		.phystatus2           (),                                                      //                    .phystatus2
		.phystatus3           (),                                                      //                    .phystatus3
		.phystatus4           (),                                                      //                    .phystatus4
		.phystatus5           (),                                                      //                    .phystatus5
		.phystatus6           (),                                                      //                    .phystatus6
		.phystatus7           (),                                                      //                    .phystatus7
		.rxdata0              (),                                                      //                    .rxdata0
		.rxdata1              (),                                                      //                    .rxdata1
		.rxdata2              (),                                                      //                    .rxdata2
		.rxdata3              (),                                                      //                    .rxdata3
		.rxdata4              (),                                                      //                    .rxdata4
		.rxdata5              (),                                                      //                    .rxdata5
		.rxdata6              (),                                                      //                    .rxdata6
		.rxdata7              (),                                                      //                    .rxdata7
		.rxdatak0             (),                                                      //                    .rxdatak0
		.rxdatak1             (),                                                      //                    .rxdatak1
		.rxdatak2             (),                                                      //                    .rxdatak2
		.rxdatak3             (),                                                      //                    .rxdatak3
		.rxdatak4             (),                                                      //                    .rxdatak4
		.rxdatak5             (),                                                      //                    .rxdatak5
		.rxdatak6             (),                                                      //                    .rxdatak6
		.rxdatak7             (),                                                      //                    .rxdatak7
		.rxelecidle0          (),                                                      //                    .rxelecidle0
		.rxelecidle1          (),                                                      //                    .rxelecidle1
		.rxelecidle2          (),                                                      //                    .rxelecidle2
		.rxelecidle3          (),                                                      //                    .rxelecidle3
		.rxelecidle4          (),                                                      //                    .rxelecidle4
		.rxelecidle5          (),                                                      //                    .rxelecidle5
		.rxelecidle6          (),                                                      //                    .rxelecidle6
		.rxelecidle7          (),                                                      //                    .rxelecidle7
		.rxstatus0            (),                                                      //                    .rxstatus0
		.rxstatus1            (),                                                      //                    .rxstatus1
		.rxstatus2            (),                                                      //                    .rxstatus2
		.rxstatus3            (),                                                      //                    .rxstatus3
		.rxstatus4            (),                                                      //                    .rxstatus4
		.rxstatus5            (),                                                      //                    .rxstatus5
		.rxstatus6            (),                                                      //                    .rxstatus6
		.rxstatus7            (),                                                      //                    .rxstatus7
		.rxvalid0             (),                                                      //                    .rxvalid0
		.rxvalid1             (),                                                      //                    .rxvalid1
		.rxvalid2             (),                                                      //                    .rxvalid2
		.rxvalid3             (),                                                      //                    .rxvalid3
		.rxvalid4             (),                                                      //                    .rxvalid4
		.rxvalid5             (),                                                      //                    .rxvalid5
		.rxvalid6             (),                                                      //                    .rxvalid6
		.rxvalid7             (),                                                      //                    .rxvalid7
		.test_in              (pcie2_hip_ctrl_test_in),                                //            hip_ctrl.test_in
		.simu_mode_pipe       (pcie2_hip_ctrl_simu_mode_pipe),                         //                    .simu_mode_pipe
		.rxdataskip0          (1'b0),                                                  //         (terminated)
		.rxdataskip1          (1'b0),                                                  //         (terminated)
		.rxdataskip2          (1'b0),                                                  //         (terminated)
		.rxdataskip3          (1'b0),                                                  //         (terminated)
		.rxdataskip4          (1'b0),                                                  //         (terminated)
		.rxdataskip5          (1'b0),                                                  //         (terminated)
		.rxdataskip6          (1'b0),                                                  //         (terminated)
		.rxdataskip7          (1'b0),                                                  //         (terminated)
		.rxblkst0             (1'b0),                                                  //         (terminated)
		.rxblkst1             (1'b0),                                                  //         (terminated)
		.rxblkst2             (1'b0),                                                  //         (terminated)
		.rxblkst3             (1'b0),                                                  //         (terminated)
		.rxblkst4             (1'b0),                                                  //         (terminated)
		.rxblkst5             (1'b0),                                                  //         (terminated)
		.rxblkst6             (1'b0),                                                  //         (terminated)
		.rxblkst7             (1'b0),                                                  //         (terminated)
		.rxsynchd0            (2'b00),                                                 //         (terminated)
		.rxsynchd1            (2'b00),                                                 //         (terminated)
		.rxsynchd2            (2'b00),                                                 //         (terminated)
		.rxsynchd3            (2'b00),                                                 //         (terminated)
		.rxsynchd4            (2'b00),                                                 //         (terminated)
		.rxsynchd5            (2'b00),                                                 //         (terminated)
		.rxsynchd6            (2'b00),                                                 //         (terminated)
		.rxsynchd7            (2'b00),                                                 //         (terminated)
		.rxfreqlocked0        (1'b0),                                                  //         (terminated)
		.rxfreqlocked1        (1'b0),                                                  //         (terminated)
		.rxfreqlocked2        (1'b0),                                                  //         (terminated)
		.rxfreqlocked3        (1'b0),                                                  //         (terminated)
		.rxfreqlocked4        (1'b0),                                                  //         (terminated)
		.rxfreqlocked5        (1'b0),                                                  //         (terminated)
		.rxfreqlocked6        (1'b0),                                                  //         (terminated)
		.rxfreqlocked7        (1'b0),                                                  //         (terminated)
		.currentcoeff0        (),                                                      //         (terminated)
		.currentcoeff1        (),                                                      //         (terminated)
		.currentcoeff2        (),                                                      //         (terminated)
		.currentcoeff3        (),                                                      //         (terminated)
		.currentcoeff4        (),                                                      //         (terminated)
		.currentcoeff5        (),                                                      //         (terminated)
		.currentcoeff6        (),                                                      //         (terminated)
		.currentcoeff7        (),                                                      //         (terminated)
		.currentrxpreset0     (),                                                      //         (terminated)
		.currentrxpreset1     (),                                                      //         (terminated)
		.currentrxpreset2     (),                                                      //         (terminated)
		.currentrxpreset3     (),                                                      //         (terminated)
		.currentrxpreset4     (),                                                      //         (terminated)
		.currentrxpreset5     (),                                                      //         (terminated)
		.currentrxpreset6     (),                                                      //         (terminated)
		.currentrxpreset7     (),                                                      //         (terminated)
		.txsynchd0            (),                                                      //         (terminated)
		.txsynchd1            (),                                                      //         (terminated)
		.txsynchd2            (),                                                      //         (terminated)
		.txsynchd3            (),                                                      //         (terminated)
		.txsynchd4            (),                                                      //         (terminated)
		.txsynchd5            (),                                                      //         (terminated)
		.txsynchd6            (),                                                      //         (terminated)
		.txsynchd7            (),                                                      //         (terminated)
		.txblkst0             (),                                                      //         (terminated)
		.txblkst1             (),                                                      //         (terminated)
		.txblkst2             (),                                                      //         (terminated)
		.txblkst3             (),                                                      //         (terminated)
		.txblkst4             (),                                                      //         (terminated)
		.txblkst5             (),                                                      //         (terminated)
		.txblkst6             (),                                                      //         (terminated)
		.txblkst7             ()                                                       //         (terminated)
	);

	pcie_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pcie1_coreclkout_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	pcie_system_mm_interconnect_0 mm_interconnect_0 (
		.pcie1_coreclkout_clk                              (pcie1_coreclkout_clk),                                  //                            pcie1_coreclkout.clk
		.intel_lw_uart_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // intel_lw_uart_0_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                    //    sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.pcie1_Rxm_BAR0_address                            (pcie1_rxm_bar0_address),                                //                              pcie1_Rxm_BAR0.address
		.pcie1_Rxm_BAR0_waitrequest                        (pcie1_rxm_bar0_waitrequest),                            //                                            .waitrequest
		.pcie1_Rxm_BAR0_burstcount                         (pcie1_rxm_bar0_burstcount),                             //                                            .burstcount
		.pcie1_Rxm_BAR0_byteenable                         (pcie1_rxm_bar0_byteenable),                             //                                            .byteenable
		.pcie1_Rxm_BAR0_read                               (pcie1_rxm_bar0_read),                                   //                                            .read
		.pcie1_Rxm_BAR0_readdata                           (pcie1_rxm_bar0_readdata),                               //                                            .readdata
		.pcie1_Rxm_BAR0_readdatavalid                      (pcie1_rxm_bar0_readdatavalid),                          //                                            .readdatavalid
		.pcie1_Rxm_BAR0_write                              (pcie1_rxm_bar0_write),                                  //                                            .write
		.pcie1_Rxm_BAR0_writedata                          (pcie1_rxm_bar0_writedata),                              //                                            .writedata
		.intel_lw_uart_0_s1_address                        (mm_interconnect_0_intel_lw_uart_0_s1_address),          //                          intel_lw_uart_0_s1.address
		.intel_lw_uart_0_s1_write                          (mm_interconnect_0_intel_lw_uart_0_s1_write),            //                                            .write
		.intel_lw_uart_0_s1_read                           (mm_interconnect_0_intel_lw_uart_0_s1_read),             //                                            .read
		.intel_lw_uart_0_s1_readdata                       (mm_interconnect_0_intel_lw_uart_0_s1_readdata),         //                                            .readdata
		.intel_lw_uart_0_s1_writedata                      (mm_interconnect_0_intel_lw_uart_0_s1_writedata),        //                                            .writedata
		.sysid_qsys_0_control_slave_address                (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //                  sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata               (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)  //                                            .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~rst_125_reset_n),               // reset_in0.reset
		.clk            (clk_125_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pcie1_nreset_status_reset),         // reset_in0.reset
		.clk            (pcie1_coreclkout_clk),               //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~rst_125_reset_n),                   // reset_in0.reset
		.reset_in1      (~pcie1_nreset_status_reset),         // reset_in1.reset
		.clk            (pcie1_coreclkout_clk),               //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
