// vroom_system.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module vroom_system (
		input  wire  clk_clk,                    //             clk.clk
		input  wire  reset_reset_n,              //           reset.reset_n
		input  wire  vroom_0_uart_rx_new_signal, // vroom_0_uart_rx.new_signal
		output wire  vroom_0_uart_tx_new_signal  // vroom_0_uart_tx.new_signal
	);

	wire         pll_0_outclk0_clk;                          // pll_0:outclk_0 -> [RAM:clk, ROM:clk, VROOM_0:clk, interrupt_connections_1:clk, mm_interconnect_0:pll_0_outclk0_clk, reset_controller_0:clk, rst_controller:clk]
	wire  [63:0] interrupt_connections_1_signals_new_signal; // interrupt_connections_1:irqs -> VROOM_0:irqs
	wire         vroom_0_avalon_master_waitrequest;          // mm_interconnect_0:VROOM_0_avalon_master_waitrequest -> VROOM_0:av_waitrequest
	wire  [31:0] vroom_0_avalon_master_readdata;             // mm_interconnect_0:VROOM_0_avalon_master_readdata -> VROOM_0:av_readdata
	wire  [31:0] vroom_0_avalon_master_address;              // VROOM_0:av_address -> mm_interconnect_0:VROOM_0_avalon_master_address
	wire         vroom_0_avalon_master_read;                 // VROOM_0:av_read -> mm_interconnect_0:VROOM_0_avalon_master_read
	wire   [3:0] vroom_0_avalon_master_byteenable;           // VROOM_0:av_byteenable -> mm_interconnect_0:VROOM_0_avalon_master_byteenable
	wire         vroom_0_avalon_master_readdatavalid;        // mm_interconnect_0:VROOM_0_avalon_master_readdatavalid -> VROOM_0:av_readdatavalid
	wire   [1:0] vroom_0_avalon_master_response;             // mm_interconnect_0:VROOM_0_avalon_master_response -> VROOM_0:av_response
	wire  [31:0] vroom_0_avalon_master_writedata;            // VROOM_0:av_writedata -> mm_interconnect_0:VROOM_0_avalon_master_writedata
	wire         vroom_0_avalon_master_write;                // VROOM_0:av_write -> mm_interconnect_0:VROOM_0_avalon_master_write
	wire         vroom_0_avalon_master_writeresponsevalid;   // mm_interconnect_0:VROOM_0_avalon_master_writeresponsevalid -> VROOM_0:av_writeresponsevalid
	wire   [4:0] vroom_0_avalon_master_burstcount;           // VROOM_0:av_burstcount -> mm_interconnect_0:VROOM_0_avalon_master_burstcount
	wire         mm_interconnect_0_rom_s1_chipselect;        // mm_interconnect_0:ROM_s1_chipselect -> ROM:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;          // ROM:readdata -> mm_interconnect_0:ROM_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;       // mm_interconnect_0:ROM_s1_debugaccess -> ROM:debugaccess
	wire  [14:0] mm_interconnect_0_rom_s1_address;           // mm_interconnect_0:ROM_s1_address -> ROM:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;        // mm_interconnect_0:ROM_s1_byteenable -> ROM:byteenable
	wire         mm_interconnect_0_rom_s1_write;             // mm_interconnect_0:ROM_s1_write -> ROM:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;         // mm_interconnect_0:ROM_s1_writedata -> ROM:writedata
	wire         mm_interconnect_0_rom_s1_clken;             // mm_interconnect_0:ROM_s1_clken -> ROM:clken
	wire         mm_interconnect_0_ram_s1_chipselect;        // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;          // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [12:0] mm_interconnect_0_ram_s1_address;           // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;        // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;             // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;         // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;             // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         rst_controller_reset_out_reset;             // rst_controller:reset_out -> [RAM:reset, ROM:reset, VROOM_0:rst, mm_interconnect_0:VROOM_0_reset_sink_reset_bridge_in_reset_reset]
	wire         rst_controller_reset_out_reset_req;         // rst_controller:reset_req -> [RAM:reset_req, ROM:reset_req, rst_translator:reset_req_in]
	wire         reset_controller_0_reset_out_reset;         // reset_controller_0:reset_out -> rst_controller:reset_in0

	vroom_system_RAM ram (
		.clk        (pll_0_outclk0_clk),                   //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	vroom_system_ROM rom (
		.clk         (pll_0_outclk0_clk),                    //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	CoreWrapper #(
		.SIMULATION (0)
	) vroom_0 (
		.clk                   (pll_0_outclk0_clk),                          //         clock.clk
		.av_waitrequest        (vroom_0_avalon_master_waitrequest),          // avalon_master.waitrequest
		.av_readdata           (vroom_0_avalon_master_readdata),             //              .readdata
		.av_readdatavalid      (vroom_0_avalon_master_readdatavalid),        //              .readdatavalid
		.av_response           (vroom_0_avalon_master_response),             //              .response
		.av_writeresponsevalid (vroom_0_avalon_master_writeresponsevalid),   //              .writeresponsevalid
		.av_burstcount         (vroom_0_avalon_master_burstcount),           //              .burstcount
		.av_writedata          (vroom_0_avalon_master_writedata),            //              .writedata
		.av_address            (vroom_0_avalon_master_address),              //              .address
		.av_write              (vroom_0_avalon_master_write),                //              .write
		.av_read               (vroom_0_avalon_master_read),                 //              .read
		.av_byteenable         (vroom_0_avalon_master_byteenable),           //              .byteenable
		.rst                   (rst_controller_reset_out_reset),             //    reset_sink.reset
		.irqs                  (interrupt_connections_1_signals_new_signal), //    interrupts.new_signal
		.uart_rx               (vroom_0_uart_rx_new_signal),                 //       uart_rx.new_signal
		.uart_tx               (vroom_0_uart_tx_new_signal)                  //       uart_tx.new_signal
	);

	interrupt_connections interrupt_connections_1 (
		.irqs (interrupt_connections_1_signals_new_signal), // signals.new_signal
		.clk  (pll_0_outclk0_clk)                           //   clock.clk
	);

	vroom_system_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_0 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (reset_controller_0_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	vroom_system_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                              (pll_0_outclk0_clk),                        //                            pll_0_outclk0.clk
		.VROOM_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),           // VROOM_0_reset_sink_reset_bridge_in_reset.reset
		.VROOM_0_avalon_master_address                  (vroom_0_avalon_master_address),            //                    VROOM_0_avalon_master.address
		.VROOM_0_avalon_master_waitrequest              (vroom_0_avalon_master_waitrequest),        //                                         .waitrequest
		.VROOM_0_avalon_master_burstcount               (vroom_0_avalon_master_burstcount),         //                                         .burstcount
		.VROOM_0_avalon_master_byteenable               (vroom_0_avalon_master_byteenable),         //                                         .byteenable
		.VROOM_0_avalon_master_read                     (vroom_0_avalon_master_read),               //                                         .read
		.VROOM_0_avalon_master_readdata                 (vroom_0_avalon_master_readdata),           //                                         .readdata
		.VROOM_0_avalon_master_readdatavalid            (vroom_0_avalon_master_readdatavalid),      //                                         .readdatavalid
		.VROOM_0_avalon_master_write                    (vroom_0_avalon_master_write),              //                                         .write
		.VROOM_0_avalon_master_writedata                (vroom_0_avalon_master_writedata),          //                                         .writedata
		.VROOM_0_avalon_master_response                 (vroom_0_avalon_master_response),           //                                         .response
		.VROOM_0_avalon_master_writeresponsevalid       (vroom_0_avalon_master_writeresponsevalid), //                                         .writeresponsevalid
		.RAM_s1_address                                 (mm_interconnect_0_ram_s1_address),         //                                   RAM_s1.address
		.RAM_s1_write                                   (mm_interconnect_0_ram_s1_write),           //                                         .write
		.RAM_s1_readdata                                (mm_interconnect_0_ram_s1_readdata),        //                                         .readdata
		.RAM_s1_writedata                               (mm_interconnect_0_ram_s1_writedata),       //                                         .writedata
		.RAM_s1_byteenable                              (mm_interconnect_0_ram_s1_byteenable),      //                                         .byteenable
		.RAM_s1_chipselect                              (mm_interconnect_0_ram_s1_chipselect),      //                                         .chipselect
		.RAM_s1_clken                                   (mm_interconnect_0_ram_s1_clken),           //                                         .clken
		.ROM_s1_address                                 (mm_interconnect_0_rom_s1_address),         //                                   ROM_s1.address
		.ROM_s1_write                                   (mm_interconnect_0_rom_s1_write),           //                                         .write
		.ROM_s1_readdata                                (mm_interconnect_0_rom_s1_readdata),        //                                         .readdata
		.ROM_s1_writedata                               (mm_interconnect_0_rom_s1_writedata),       //                                         .writedata
		.ROM_s1_byteenable                              (mm_interconnect_0_rom_s1_byteenable),      //                                         .byteenable
		.ROM_s1_chipselect                              (mm_interconnect_0_rom_s1_chipselect),      //                                         .chipselect
		.ROM_s1_clken                                   (mm_interconnect_0_rom_s1_clken),           //                                         .clken
		.ROM_s1_debugaccess                             (mm_interconnect_0_rom_s1_debugaccess)      //                                         .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_controller_0_reset_out_reset), // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
