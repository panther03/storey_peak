
module vroom_system (
	clk_clk,
	reset_reset_n,
	vroom_0_uart_rx_new_signal,
	vroom_0_uart_tx_new_signal);	

	input		clk_clk;
	input		reset_reset_n;
	input		vroom_0_uart_rx_new_signal;
	output		vroom_0_uart_tx_new_signal;
endmodule
