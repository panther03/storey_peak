// jtag_uart.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module jtag_uart (
		input  wire        av_chipselect,  //    av.chipselect
		input  wire        av_address,     //      .address
		input  wire        av_read_n,      //      .read_n
		output wire [31:0] av_readdata,    //      .readdata
		input  wire        av_write_n,     //      .write_n
		input  wire [31:0] av_writedata,   //      .writedata
		output wire        av_waitrequest, //      .waitrequest
		input  wire        clk_clk,        //   clk.clk
		output wire        irq_irq,        //   irq.irq
		input  wire        reset_reset_n   // reset.reset_n
	);

	jtag_uart_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),        //               clk.clk
		.rst_n          (reset_reset_n),  //             reset.reset_n
		.av_chipselect  (av_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (av_address),     //                  .address
		.av_read_n      (av_read_n),      //                  .read_n
		.av_readdata    (av_readdata),    //                  .readdata
		.av_write_n     (av_write_n),     //                  .write_n
		.av_writedata   (av_writedata),   //                  .writedata
		.av_waitrequest (av_waitrequest), //                  .waitrequest
		.av_irq         (irq_irq)         //               irq.irq
	);

endmodule
